module score_rom ( input [8:0]	addr,
						output [15:0]	data
					 );
	parameter ADDR_WIDTH = 9;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;			
	// ROM definition				
	parameter [0:239][15:0] ROM = {
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000111111111000,   
	16'b0001111111111000,   
	16'b0001100000000000,  
	16'b0001100000000000,   
	16'b0001111111111000,   
	16'b0000111111111000,   
	16'b0000000000011000,   
	16'b0000000000011000,   
	16'b0001111111111000,   
	16'b0001111111110000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000, 

	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000111111111000,   
	16'b0001111111111000,   
	16'b0001100000000000,   
	16'b0001100000000000,   
	16'b0001100000000000,   
	16'b0001100000000000,   
	16'b0001100000000000,   
	16'b0001100000000000,   
	16'b0001111111111000,   
	16'b0000111111111000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000, 

	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000111111110000,   
	16'b0001111111111000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001111111111000,   
	16'b0000111111110000,   
	16'b0000000000000000,
	16'b0000000000000000,   
	16'b0000000000000000,

	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000111111110000,   
	16'b0001111111111000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001111111111000,   
	16'b0001111111110000,   
	16'b0001100111000000,   
	16'b0001100011100000,   
	16'b0001100001110000,   
	16'b0001100000111000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,

	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0001111111111000,   
	16'b0001111111111000,   
	16'b0001100000000000,   
	16'b0001100000000000,   
	16'b0001111111111000,   
	16'b0001111111111000,   
	16'b0001100000000000,   
	16'b0001100000000000,   
	16'b0001111111111000,   
	16'b0001111111111000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000, 

	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000111111110000,   
	16'b0001111111111000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001100000011000,   
	16'b0001111111111000,   
	16'b0000111111110000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,

	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000001111000000,   
	16'b0000011111000000,   
	16'b0000111111000000,   
	16'b0000000111000000,   
	16'b0000000111000000,   
	16'b0000000111000000,   
	16'b0000000111000000,   
	16'b0000000111000000,   
	16'b0000000111000000,   
	16'b0000000111000000,   
	16'b0000000000000000,   
	16'b0000000000000000,   
	16'b0000000000000000, 

	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000111111110000,  
	16'b0001111111111000,  
	16'b0001110000111000,  
	16'b0000000000111000,  
	16'b0000000001110000,  
	16'b0000000011100000,  
	16'b0000000111000000,  
	16'b0000001110000000,  
	16'b0000111111111000,  
	16'b0001111111111000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,

	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000111111110000,  
	16'b0001111111111000,  
	16'b0001100000011000,  
	16'b0000000000011000,  
	16'b0000000111110000,  
	16'b0000000111110000,  
	16'b0000000000011000,  
	16'b0001100000011000,  
	16'b0001111111111000,  
	16'b0000111111110000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,

	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000011111000,  
	16'b0000000111111000,  
	16'b0000001110011000,  
	16'b0000011100011000,  
	16'b0000111000011000,  
	16'b0001111111111100,  
	16'b0001111111111100,  
	16'b0000000000011000,  
	16'b0000000000011000,  
	16'b0000000000011000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,

	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0001111111111000,  
	16'b0001111111111000,  
	16'b0001100000000000,  
	16'b0001100000000000,  
	16'b0001111111110000,  
	16'b0001111111111000,  
	16'b0000000000011000,  
	16'b0001100000011000,  
	16'b0001111111111000,  
	16'b0000111111110000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,

	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000111111110000,  
	16'b0001111111111000,  
	16'b0001100000011000,  
	16'b0001100000000000,  
	16'b0001111111110000,  
	16'b0001111111111000,  
	16'b0001100000011000,  
	16'b0001100000011000,  
	16'b0001111111111000, 
	16'b0000111111110000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,

	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0001111111111000,  
	16'b0001111111111000,  
	16'b0000000001110000,  
	16'b0000000001110000,  
	16'b0000000011100000,  
	16'b0000000011100000,  
	16'b0000000111000000,  
	16'b0000000111000000,  
	16'b0000001110000000,  
	16'b0000001110000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,

	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000111111110000,  
	16'b0001111111111000,  
	16'b0001100000011000,  
	16'b0001100000011000,  
	16'b0000111111110000,  
	16'b0000111111110000,  
	16'b0001100000011000,  
	16'b0001100000011000,  
	16'b0001111111111000,  
	16'b0000111111110000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,

	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000111111110000,  
	16'b0001111111111000,  
	16'b0001100000011000,  
	16'b0001100000011000,  
	16'b0001111111111000,  
	16'b0000111111111000,  
	16'b0000000000011000,  
	16'b0001100000011000,  
	16'b0001111111111000,  
	16'b0000111111110000,  
	16'b0000000000000000,  
	16'b0000000000000000,  
	16'b0000000000000000,
	};
	assign data = ROM[addr];
endmodule