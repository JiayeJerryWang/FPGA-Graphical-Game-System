module pac_rom ( input [6:0]	addr,
						output [15:0]	data
					 );

	parameter ADDR_WIDTH = 7;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:95][DATA_WIDTH-1:0] ROM = {
			16'b0000011111110000, // left x01
			16'b0000111111111000,
			16'b0001111111111100,
			16'b0011111111111111,
			16'b0011111111111110,
			16'b0111111111111100,
			16'b0111111111111000,
			16'b0111111111100000,
			16'b0111111111100000,
			16'b0011111111111000,
			16'b0011111111111100,
			16'b0011111111111110,
			16'b0011111111111111,
			16'b0001111111111100,
			16'b0000111111111000,
			16'b0000011111110000,
		  
         
			16'b0000111111110000, // closed x02
			16'b0001111111111000,
			16'b0011111111111100,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0111111111111110,
			16'b0011111111111100,
			16'b0001111111111000,
			16'b0000111111110000,

			16'b0000111111110000,
			16'b0011111111111100,
			16'b1110011111100111,
			16'b1101101111011011,
			16'b1110011111100111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111001111100111,
			16'b1110000111000011,
			16'b1100000010000001,
		  
			16'b0001000000001000, //up x04
			16'b0001100000011000,
			16'b0011110000111100,
			16'b0111111001111110,
			16'b1111111001111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b0111111111111110,
			16'b0011111111111100,
			16'b0001111111111000,
			16'b0000000110000000,
			16'b0000000000000000,

			16'b0000000000000000, // down x05
			16'b0000000110000000,
			16'b0001111111111000,
			16'b0011111111111100,
			16'b0111111111111110,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111111111111,
			16'b1111111001111111,
			16'b0111111001111110,
			16'b0011110000111100,
			16'b0001100000011000,
			16'b0001000000001000,

			16'b0000111111100000, // right x06
			16'b0001111111110000,
			16'b0011111111111000,
			16'b1111111111111100,
			16'b0111111111111100,
			16'b0011111111111110,
			16'b0001111111111110,
			16'b0000011111111110,
			16'b0000011111111110,
			16'b0001111111111110,
			16'b0011111111111100,
			16'b0111111111111100,
			16'b1111111111111100,
			16'b0011111111111000,
			16'b0001111111110000,
			16'b0000111111100000
			};

	assign data = ROM[addr];

endmodule  
//module pac_rom ( input [5:0]	addr,
//						output [26:0]	data
//					 );
//
//	parameter ADDR_WIDTH = 16;
//   parameter DATA_WIDTH =  16;
//	logic [ADDR_WIDTH-1:0] addr_reg;
//	// ROM definition
//	parameter [0:ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
//	16'b0000000000000000,  
//	16'b0000011111100000,
//	16'b0001111111111000,
//	16'b0011111111111100,
//	16'b0111111111111110,
//	16'b1111111111111110,
//	16'b1111111111100000,
//	16'b1111111000000000,
//	16'b1111111000000000,
//	16'b1111111111100000,
//	16'b1111111111111110,
//	16'b0111111111111110,
//	16'b0011111111111100,
//	16'b0001111111111000,
//	16'b0000011111100000,
//	16'b0000000000000000
//	};
//
//	assign data = ROM[addr];
//
//endmodule

// 
// sprite_dot_small( 0) <= "0000000000000000";
// sprite_dot_small( 1) <= "0000000000000000";
// sprite_dot_small( 2) <= "0000000000000000";
// sprite_dot_small( 3) <= "0000000000000000";
// sprite_dot_small( 4) <= "0000000000000000";
// sprite_dot_small( 5) <= "0000000000000000";
// sprite_dot_small( 6) <= "0000000110000000";
// sprite_dot_small( 7) <= "0000001111000000";
// sprite_dot_small( 8) <= "0000000110000000";
// sprite_dot_small( 9) <= "0000000000000000";
// sprite_dot_small(10) <= "0000000000000000";
// sprite_dot_small(11) <= "0000000000000000";
// sprite_dot_small(12) <= "0000000000000000";
// sprite_dot_small(13) <= "0000000000000000";
// sprite_dot_small(14) <= "0000000000000000";
// sprite_dot_small(15) <= "0000000000000000";
// 
// sprite_dot_large( 0) <= "0000000000000000";
// sprite_dot_large( 1) <= "0000000000000000";
// sprite_dot_large( 2) <= "0000000000000000";
// sprite_dot_large( 3) <= "0000001111000000";
// sprite_dot_large( 4) <= "0000011111100000";
// sprite_dot_large( 5) <= "0000111111110000";
// sprite_dot_large( 6) <= "0001111111111000";
// sprite_dot_large( 7) <= "0001111111111000";
// sprite_dot_large( 8) <= "0001111111111000";
// sprite_dot_large( 9) <= "0000111111110000";
// sprite_dot_large(10) <= "0000011111100000";
// sprite_dot_large(11) <= "0000001111000000";
// sprite_dot_large(12) <= "0000000000000000";
// sprite_dot_large(13) <= "0000000000000000";
// sprite_dot_large(14) <= "0000000000000000";
// sprite_dot_large(15) <= "0000000000000000"; 
// 
// sprite_ghost( 0) <= "0000000000000000";
// sprite_ghost( 1) <= "0000111111110000";
// sprite_ghost( 2) <= "0111111111111110";
// sprite_ghost( 3) <= "1111111111111111";
// sprite_ghost( 4) <= "1111111111111111";
// sprite_ghost( 5) <= "1111000111100011";
// sprite_ghost( 6) <= "1111000111100011";
// sprite_ghost( 7) <= "1111111111111111";
// sprite_ghost( 8) <= "1111111111111111";
// sprite_ghost( 9) <= "1111111111111111";
// sprite_ghost(10) <= "1111111111111111";
// sprite_ghost(11) <= "1111111111111111";
// sprite_ghost(12) <= "1111111111111111";
// sprite_ghost(13) <= "1111111111111111";
// sprite_ghost(14) <= "1101111001111011";
// sprite_ghost(15) <= "1000110000110001"; 


//
//module spriteData ( input [7:0]	addr,
//						output [31:0]	data
//					 );
//
//	parameter ADDR_WIDTH = 8;
//   parameter DATA_WIDTH =  32;
//	logic [ADDR_WIDTH-1:0] addr_reg;
//
//	// ROM definition
//	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
//
//		//Pacman facing left
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000001111111000000000000,
//		32'b 00000000000111111111111000000000,
//		32'b 00000000011111111111111110000000,
//		32'b 00000000111111111111111111000000,
//		32'b 00000011111111111111111111100000,
//		32'b 00000111111111111111111110000000,
//		32'b 00001111111111111111111000000000,
//		32'b 00001111111111111111110000000000,
//		32'b 00001111111111111111000000000000,
//		32'b 00011111111111111000000000000000,
//		32'b 00011111111111110000000000000000,
//		32'b 00011111111111111000000000000000,
//		32'b 00001111111111111111000000000000,
//		32'b 00001111111111111111110000000000,
//		32'b 00001111111111111111111000000000,
//		32'b 00000111111111111111111110000000,
//		32'b 00000011111111111111111111100000,
//		32'b 00000000111111111111111111000000,
//		32'b 00000000011111111111111110000000,
//		32'b 00000000000111111111111000000000,
//		32'b 00000000000001111111000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//
//		//Pacman facing left
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000011111110000000000000,
//		32'b 00000000011111111111100000000000,
//		32'b 00000001111111111111111000000000,
//		32'b 00000011111111111111111100000000,
//		32'b 00000111111111111111111111000000,
//		32'b 00000001111111111111111111100000,
//		32'b 00000000011111111111111111110000,
//		32'b 00000000001111111111111111110000,
//		32'b 00000000000011111111111111110000,
//		32'b 00000000000000011111111111111000,
//		32'b 00000000000000001111111111111000,
//		32'b 00000000000000011111111111111000,
//		32'b 00000000000011111111111111110000,
//		32'b 00000000001111111111111111110000,
//		32'b 00000000011111111111111111110000,
//		32'b 00000001111111111111111111100000,
//		32'b 00000111111111111111111111000000,
//		32'b 00000011111111111111111100000000,
//		32'b 00000001111111111111111000000000,
//		32'b 00000000011111111111100000000000,
//		32'b 00000000000011111110000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//
//		//Pacman facing up
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000100000000001000000000,
//		32'b 00000000011100000000001110000000,
//		32'b 00000000111100000000001111000000,
//		32'b 00000011111100000000001111100000,
//		32'b 00000111111110000000011111100000,
//		32'b 00001111111110000000011111110000,
//		32'b 00001111111111000000111111110000,
//		32'b 00001111111111000000111111110000,
//		32'b 00011111111111100001111111110000,
//		32'b 00011111111111100011111111110000,
//		32'b 00011111111111110111111111111000,
//		32'b 00001111111111111111111111110000,
//		32'b 00001111111111111111111111110000,
//		32'b 00001111111111111111111111110000,
//		32'b 00000111111111111111111111100000,
//		32'b 00000011111111111111111111100000,
//		32'b 00000000111111111111111111000000,
//		32'b 00000000011111111111111110000000,
//		32'b 00000000000111111111111000000000,
//		32'b 00000000000001111111000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//
//		//Pacman facing down
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000001111111000000000000,
//		32'b 00000000000111111111111000000000,
//		32'b 00000000011111111111111110000000,
//		32'b 00000000111111111111111111000000,
//		32'b 00000011111111111111111111100000,
//		32'b 00000111111111111111111111100000,
//		32'b 00001111111111111111111111110000,
//		32'b 00001111111111111111111111110000,
//		32'b 00001111111111111111111111110000,
//		32'b 00011111111111111011111111111000,
//		32'b 00011111111111110001111111111000,
//		32'b 00011111111111100001111111111000,
//		32'b 00001111111111000000111111110000,
//		32'b 00001111111111000000111111110000,
//		32'b 00001111111110000000011111110000,
//		32'b 00000111111110000000011111100000,
//		32'b 00000011111100000000001111100000,
//		32'b 00000000111100000000001111000000,
//		32'b 00000000011100000000001110000000,
//		32'b 00000000000100000000001000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//
//		//Ghost sprite
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000111111111110000000000,
//		32'b 00000000011111111111111000000000,
//		32'b 00000000111111111111111100000000,
//		32'b 00000001111111111111111110000000,
//		32'b 00000011111111111111111111000000,
//		32'b 00000111111111111111111111100000,
//		32'b 00000111110011111111100111100000,
//		32'b 00001111100001111111000011110000,
//		32'b 00001111100001111111000011110000,
//		32'b 00001111100001111111000011110000,
//		32'b 00011111110011111111100111111000,
//		32'b 00011111111111111111111111111000,
//		32'b 00011111111111111111111111111000,
//		32'b 00011111111111111111111111111000,
//		32'b 00011111111111111111111111111000,
//		32'b 00011111111111111111111111111000,
//		32'b 00011110111111110111111110111000,
//		32'b 00011100011111100011111100011000,
//		32'b 00011100001111100001111000011000,
//		32'b 00011000000111000000111000011000,
//		32'b 00010000000010000000010000001000,
//		32'b 00010000000010000000010000001000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000,
//		32'b 00000000000000000000000000000000
//
//	};
//
//	assign data = ROM[addr];
//
//endmodule