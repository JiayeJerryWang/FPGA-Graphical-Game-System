module dot_rom ( input [5:0]	addr,
						output [15:0]	data
					 );

	parameter ADDR_WIDTH = 7;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;			
	// ROM definition				
	parameter [0:15][15:0] ROM = {
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000110000000,
	16'b0000001111000000,
	16'b0000000110000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000,
	16'b0000000000000000
	};

	assign data = ROM[addr];
endmodule



