module start_rom ( input [5:0]	addr,
						output [39:0]	data
					 );
	parameter ADDR_WIDTH = 6;
   parameter DATA_WIDTH =  40;
	logic [ADDR_WIDTH-1:0] addr_reg;
	parameter [0:29][39:0] rom = {
  40'b0000000000000000000000000000000000000000,         
  40'b0000000000000000000000000000000000000000, 
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,  
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0111110011111110000100000011111001111111,
  40'b1000000000010000001010000010001000001000,
  40'b0111100000010000010001000011111000001000,
  40'b0000010000010000111111100011000000001000,
  40'b0000010000010001000000010010100000001000,
  40'b1111100000010001000000010010001100001000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
  40'b0000000000000000000000000000000000000000,
		};
		assign data = rom[addr];
endmodule