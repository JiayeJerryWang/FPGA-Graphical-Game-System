module died_rom ( input [5:0]	addr,
						output [39:0]	data
					 );
	parameter ADDR_WIDTH = 6;
   parameter DATA_WIDTH =  40;
	logic [ADDR_WIDTH-1:0] addr_reg;
	parameter [0:29][39:0] rom = {
		40'b0000000000000000000000000000000000000000,         
		40'b0000000000000000000000000000000000000000, 
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,  
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000010001001111001001000000000000000,
		40'b0000000001010001001001001000000000000000,
		40'b0000000000100001001001001000000000000000,
		40'b0000000000100001001001001000000000000000,
		40'b0000000000100001001001001000000000000000,
		40'b0000000000100001111001111000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000010000001111000011111001111111000000,
		40'b0000010000001001000100000000001000000000,
		40'b0000010000001001000011110000001000000000,
		40'b0000010000001001000000001000001000000000,
		40'b0000010000001001000000001000001000000000,
		40'b0000011111101111000111110000001000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		};
		assign data = rom[addr];
endmodule